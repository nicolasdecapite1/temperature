// module real_div(input real a, input real b, output real c);
//     initial begin
//         c <= a/b;
//     end
    
// endmodule